module shield_FSM();
endmodule