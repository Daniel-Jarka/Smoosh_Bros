module hit_FSM();
endmodule