module knockback (

);

endmodule