module ledge_FSM ();
endmodule