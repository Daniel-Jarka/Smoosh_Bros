module movement_FSM();
endmodule