module dodge_FSM ();
endmodule